module im (
  input clk,
  input [31:0] addr,
  output [31:0] data
);
  reg [31:0] mem [0:255];  
  integer i=0;
 initial begin
	for (i=0; i<250; i=i+1) mem[i] = 32'b0;//mem[i] = 32'b0; 8 addi $t0, $0, 7
    mem[40] = 32'b001000_00000_01000_0000000000000111; //addi $t0, $0, 7
	 mem[41] = 32'b001000_00000_01001_0000000000001000; //addi $t1, $0, 8
	 //mem[3] = 32'b000100_01000_01001_0000000000000001;//beq $t0, $t1, 1
	 
	 mem[42] = 32'b000011_00000_00000_0000000000001011;//jal 10;
	 mem[43] = 32'b000000_01000_01001_01010_00000_100000;//add $t2, $t0, $t1
	 mem[44] = 32'b101011_00000_01010_0000000000000000;//sw $t2, 0($t0)
	 mem[45] = 32'b000000_01000_01010_01010_00000_100000;//add $t2, $t0, $t2
	 mem[46] = 32'b100011_00000_01011_0000000000000000;//lw $t3, 0($t0)
	 mem[47] = 32'b000010_00000_00000_0000000000001101;//j 13;
	 
	 mem[12] = 32'b000000_11111_00000_00000_00000_001000; //jr $ra;
	 /*mem[2] = 32'b001000_01000_01000_0000000000000111; //addi $t0, $t0, 7
	 mem[3] = 32'b001000_00000_01001_0000000000000001; //addi $t1, $0, 1
	 mem[4] = 32'b000000_01000_01001_01010_00000_100000;//add $t2, $t0, $t1
	 mem[5] = 32'b101011_00000_01010_0000000000000000;//sw $t2, 0($t0)
	 mem[6] = 32'b100011_00000_01011_0000000000000000;//lw $t3, 0($t0)*/
	 /*mem[2] =32'h21280009;//addi $t0, $t1, 9
    mem[3] =32'h01098824;//and $s1, $t0, $t1
    mem[4] =32'h01099025;//or $s2, $t0, $t1

    mem[5] =32'hac090000;//sw $t1, 0($0)
    mem[6] =32'h8c170000;//lw $t0, 0($)
*/
    /*
    mem[1] =32'h21300010; //addi $s0, $t1, 2
mem[2]=32'h360b0000; //ori  $t3, $s0, 0
mem[3]=32'h320b0006; //andi $t3, $s0, 6
mem[4]=32'had700000; //sw   $s0, 0($t3)
mem[5]=32'h8d6c0000; //lw   $t4, 0($t3)*/

//mem[10] = 32'b001000_00000_01000_0000000000000111;
/*
  mem[1] = 32'h21480005; //   addi $t0, $t2, 5
mem[2] = 32'h0C000004; //   jal b
mem[3] = 32'h21480004; //   addi $t0, $t2, 4
mem[4] = 32'h21300002; //b: addi $s0, $t1, 2
//0000 0011 1110 0000 0000 0000 0000 1000
mem[5] = 32'h03E00008; // jr $ra
mem[6] = 32'b
*/
  end
  assign data = mem[addr>>2];
 
endmodule

